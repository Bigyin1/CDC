class packet;
        logic [64-1:0] tdata;
        logic                   tid;
endclass
